// PRCO Register Set

`include "inc/prco_constants.v"

module prco_regs (
    input               i_clk,
    input               i_en,
    input               i_reset,
    
    // Pipeline control
    input               i_p_cp,
    output reg          q_p_cp,

    input               i_p_stalled,
    input               i_p_valid,
    output              q_p_stalled,
    output reg          q_p_valid,
    input               i_p_ce,
    output              q_p_ce,

    // Dual port memory access
    input [2:0]         i_sela,
    output reg [15:0]   q_data,
    input [2:0]         i_selb,
    output reg [15:0]   q_datb,

    // Write enable pin
    input               i_we,
    input [2:0]         i_seld,
    input [15:0]        i_datd
);
    // 8 16-bit registers
    reg [15:0] r_regs[0:7]/*verilator public_flat*/;

    reg [7:0] foo /*verilator public_flat*/;
    
    // Reset interator
    integer i;

    always @(posedge i_clk, posedge i_reset, posedge i_en)
    begin
        if(i_en == 1 && q_p_ce) begin
            // Reset the register set
            if(i_reset == 1) begin
                $display("Resetting Registers");
                for(i = 0; i < 6; i = i + 1) begin
                    r_regs[i] <= 16'h0;
                end
                r_regs[`REG_SP] <= 16'h00FF;
                r_regs[`REG_BP] <= 16'h00FF;

                // Output something so we don't latch
                q_data <= 16'h0;
                q_datb <= 16'h0;
            end 
            // Return values
            else begin
                // Write to a register
                if(i_we == 1) begin
                    $display("Writing register %d value: %h",
                        i_seld, i_datd);
                    r_regs[i_seld] <= i_datd;
                end

                // Writeking output
                q_data <= r_regs[i_sela];
                q_datb <= r_regs[i_selb];
            end
        end
    end

    // Pipeline control
    // We are stalled if we are ready but the next stage isn't ready (stalled)
    assign q_p_stalled = q_p_valid && i_p_stalled;

    // Ready to progress if: previous stage is ready (valid)
    // and next stage isn't stalled.
    assign q_p_ce       = i_p_valid && !q_p_stalled;

    always @(posedge i_clk) begin
        if (q_p_stalled) begin
            $display("REG: Stalled because of dec!");
        end

        if (q_p_ce) begin
            $display("REG: doing...");
            q_p_cp <= 1;
        end else begin
            q_p_cp <= 0;
        end
    end
    
    always @(posedge i_clk) begin
        if (i_reset || i_p_cp) begin
            q_p_valid <= 0;
        end else if (q_p_ce) begin
            q_p_valid <= i_p_valid;
        end else if (i_p_ce) begin
            q_p_valid <= 0;
        end
    end

endmodule